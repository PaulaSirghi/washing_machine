library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity timer_mux is
	port(SEL2:in STD_LOGIC_VECTOR(3 downto 0);
	TIMP:out STD_LOGIC_VECTOR(15 DOWNTO 0));
end timer_mux;
architecture mux2 of timer_mux is
begin
	with SEL2 select
	TIMP <= "0000000001001001" WHEN "0000",
	"0000000001100011" WHEN "0001",
	"0000000001100100" WHEN "0010",
	"0000000001111000" WHEN "0011",
	"0000000001010000" WHEN "0100",
	"0000000001100100" WHEN "0101",
	"0000000001100110" WHEN "0110",
	"0000000010000000" WHEN "0111",
	"0000000001010001" WHEN "1000",
	"0000000001100101" WHEN "1001",
	"0000000001101000" WHEN "1010",
	"0000000010000010" WHEN "1011",
	"0000000001010010" WHEN "1100",
	"0000000001100110" WHEN "1101",
	"0000000001110000" WHEN "1110",
	"0000000010000100" WHEN others;
	
END mux2;
